virtual class Transaction;

endclass