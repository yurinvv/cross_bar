`timescale 1ns/1ns

module tb;
	
	import tb_pckg::*;
	
	/////////////////////////////////////
	//  Select the Test
	/////////////////////////////////////
	//Test0 test;
	//Test1 test;
	//Test2 test;
	//Test3 test;
	//Test4 test;
	//Test5 test;
	//Test6 test;
	//Test7 test;
	////////////////////////////////////
	
	localparam CLOCK_PERIOD = 10;

	bit aclk;
	bit aresetn;

endmodule