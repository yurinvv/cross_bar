package tb_pckg;
	`include "Transaction.svh"
	`include "RequestTransaction.svh"
	`include "RespDataTransaction.svh"
	`include "Driver.svh"
	`include "DriverReq.svh"
	`include "DriverResp.svh"
	`include "Sequencer.svh"
	`include "Monitor.svh"
	`include "MonitorResp.svh"
	`include "MonitorReq.svh"
	`include "Agent.svh"
	`include "Scoreboard.svh"
	`include "Environment.svh"
	`include "BaseTest.svh"
	`include "DirectWriteTest.svh"
	`include "DirectReadTest.svh"

endpackage