package tb_pckg;
//	`include "Driver.svh"
//	`include "OutData.svh"
//	`include "Monitor.svh"
//	`include "Scoreboard.svh"
//	`include "Environment.svh"
//	`include "BaseTest.svh"
//	`include "Test0.svh"
//	`include "Test1.svh"
//	`include "Test2.svh"
//	`include "Test3.svh"
//	`include "Test4.svh"
//	`include "Test5.svh"
//	`include "Test6.svh"
//	`include "Test7.svh"

endpackage