virtual class Transaction;
	
	
endclass