virtual class Monitor;
	int id;
	virtual cross_bar_if vif;
	mailbox fifo;
endclass